module sipo_tb;
